`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:42:27 03/05/2014 
// Design Name: 
// Module Name:    BusSplitter8_26 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module BusSplitter8_26(
    input [7:0] IN1,
    output [25:0] T1
    );

	assign T1 = IN1;

endmodule
