`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:25:30 03/01/2014 
// Design Name: 
// Module Name:    SubClock 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module SubClockDyn(
		input CLK,
		input [25:0] Freq,
		output OUTCLK
    );
	 
	 reg [25:0] wait1, div;
	 reg CLK_;
	 
	 assign OUTCLK = CLK_; // output clock
	 
	 // clear out variables
	 initial begin
		wait1 = 0;
		CLK_ = 0;
		div = 0;
	 end
	 
	 
	 always @(posedge CLK) begin
		// wait until clock hits half of the counted time.
		wait1 <= wait1+1; // count up 1
		
		case(Freq) // dividers >> 2
				1: div <= 25000000;
				2: div <= 12500000;
				3: div <= 8333333;
				4: div <= 6250000;
				5: div <= 5000000;
				6: div <= 4166667;
				7: div <= 3571429;
				8: div <= 3125000;
				9: div <= 2777778;
				10: div <= 2500000;
				11: div <= 2272727;
				12: div <= 2083333;
				13: div <= 1923077;
				14: div <= 1785714;
				15: div <= 1666667;
				16: div <= 1562500;
				17: div <= 1470588;
				18: div <= 1388889;
				19: div <= 1315789;
				20: div <= 1250000;
				21: div <= 1190476;
				22: div <= 1136364;
				23: div <= 1086957;
				24: div <= 1041667;
				25: div <= 1000000;
				26: div <= 961538;
				27: div <= 925926;
				28: div <= 892857;
				29: div <= 862069;
				30: div <= 833333;
				31: div <= 806452;
				32: div <= 781250;
				33: div <= 757576;
				34: div <= 735294;
				35: div <= 714286;
				36: div <= 694444;
				37: div <= 675676;
				38: div <= 657895;
				39: div <= 641026;
				40: div <= 625000;
				41: div <= 609756;
				42: div <= 595238;
				43: div <= 581395;
				44: div <= 568182;
				45: div <= 555556;
				46: div <= 543478;
				47: div <= 531915;
				48: div <= 520833;
				49: div <= 510204;
				50: div <= 500000;
				51: div <= 490196;
				52: div <= 480769;
				53: div <= 471698;
				54: div <= 462963;
				55: div <= 454545;
				56: div <= 446429;
				57: div <= 438596;
				58: div <= 431034;
				59: div <= 423729;
				60: div <= 416667;
				61: div <= 409836;
				62: div <= 403226;
				63: div <= 396825;
				64: div <= 390625;
				65: div <= 384615;
				66: div <= 378788;
				67: div <= 373134;
				68: div <= 367647;
				69: div <= 362319;
				70: div <= 357143;
				71: div <= 352113;
				72: div <= 347222;
				73: div <= 342466;
				74: div <= 337838;
				75: div <= 333333;
				76: div <= 328947;
				77: div <= 324675;
				78: div <= 320513;
				79: div <= 316456;
				80: div <= 312500;
				81: div <= 308642;
				82: div <= 304878;
				83: div <= 301205;
				84: div <= 297619;
				85: div <= 294118;
				86: div <= 290698;
				87: div <= 287356;
				88: div <= 284091;
				89: div <= 280899;
				90: div <= 277778;
				91: div <= 274725;
				92: div <= 271739;
				93: div <= 268817;
				94: div <= 265957;
				95: div <= 263158;
				96: div <= 260417;
				97: div <= 257732;
				98: div <= 255102;
				99: div <= 252525;
				100: div <= 250000;
				101: div <= 247525;
				102: div <= 245098;
				103: div <= 242718;
				104: div <= 240385;
				105: div <= 238095;
				106: div <= 235849;
				107: div <= 233645;
				108: div <= 231481;
				109: div <= 229358;
				110: div <= 227273;
				111: div <= 225225;
				112: div <= 223214;
				113: div <= 221239;
				114: div <= 219298;
				115: div <= 217391;
				116: div <= 215517;
				117: div <= 213675;
				118: div <= 211864;
				119: div <= 210084;
				120: div <= 208333;
				121: div <= 206612;
				122: div <= 204918;
				123: div <= 203252;
				124: div <= 201613;
				125: div <= 200000;
				126: div <= 198413;
				127: div <= 196850;
				128: div <= 195313;
				129: div <= 193798;
				130: div <= 192308;
				131: div <= 190840;
				132: div <= 189394;
				133: div <= 187970;
				134: div <= 186567;
				135: div <= 185185;
				136: div <= 183824;
				137: div <= 182482;
				138: div <= 181159;
				139: div <= 179856;
				140: div <= 178571;
				141: div <= 177305;
				142: div <= 176056;
				143: div <= 174825;
				144: div <= 173611;
				145: div <= 172414;
				146: div <= 171233;
				147: div <= 170068;
				148: div <= 168919;
				149: div <= 167785;
				150: div <= 166667;
				151: div <= 165563;
				152: div <= 164474;
				153: div <= 163399;
				154: div <= 162338;
				155: div <= 161290;
				156: div <= 160256;
				157: div <= 159236;
				158: div <= 158228;
				159: div <= 157233;
				160: div <= 156250;
				161: div <= 155280;
				162: div <= 154321;
				163: div <= 153374;
				164: div <= 152439;
				165: div <= 151515;
				166: div <= 150602;
				167: div <= 149701;
				168: div <= 148810;
				169: div <= 147929;
				170: div <= 147059;
				171: div <= 146199;
				172: div <= 145349;
				173: div <= 144509;
				174: div <= 143678;
				175: div <= 142857;
				176: div <= 142045;
				177: div <= 141243;
				178: div <= 140449;
				179: div <= 139665;
				180: div <= 138889;
				181: div <= 138122;
				182: div <= 137363;
				183: div <= 136612;
				184: div <= 135870;
				185: div <= 135135;
				186: div <= 134409;
				187: div <= 133690;
				188: div <= 132979;
				189: div <= 132275;
				190: div <= 131579;
				191: div <= 130890;
				192: div <= 130208;
				193: div <= 129534;
				194: div <= 128866;
				195: div <= 128205;
				196: div <= 127551;
				197: div <= 126904;
				198: div <= 126263;
				199: div <= 125628;
				200: div <= 125000;
				201: div <= 124378;
				202: div <= 123762;
				203: div <= 123153;
				204: div <= 122549;
				205: div <= 121951;
				206: div <= 121359;
				207: div <= 120773;
				208: div <= 120192;
				209: div <= 119617;
				210: div <= 119048;
				211: div <= 118483;
				212: div <= 117925;
				213: div <= 117371;
				214: div <= 116822;
				215: div <= 116279;
				216: div <= 115741;
				217: div <= 115207;
				218: div <= 114679;
				219: div <= 114155;
				220: div <= 113636;
				221: div <= 113122;
				222: div <= 112613;
				223: div <= 112108;
				224: div <= 111607;
				225: div <= 111111;
				226: div <= 110619;
				227: div <= 110132;
				228: div <= 109649;
				229: div <= 109170;
				230: div <= 108696;
				231: div <= 108225;
				232: div <= 107759;
				233: div <= 107296;
				234: div <= 106838;
				235: div <= 106383;
				236: div <= 105932;
				237: div <= 105485;
				238: div <= 105042;
				239: div <= 104603;
				240: div <= 104167;
				241: div <= 103734;
				242: div <= 103306;
				243: div <= 102881;
				244: div <= 102459;
				245: div <= 102041;
				246: div <= 101626;
				247: div <= 101215;
				248: div <= 100806;
				249: div <= 100402;
				250: div <= 100000;
				251: div <= 99602;
				252: div <= 99206;
				253: div <= 98814;
				254: div <= 98425;
				255: div <= 98039;
				256: div <= 97656;
				257: div <= 97276;
				258: div <= 96899;
				259: div <= 96525;
				260: div <= 96154;
				261: div <= 95785;
				262: div <= 95420;
				263: div <= 95057;
				264: div <= 94697;
				265: div <= 94340;
				266: div <= 93985;
				267: div <= 93633;
				268: div <= 93284;
				269: div <= 92937;
				270: div <= 92593;
				271: div <= 92251;
				272: div <= 91912;
				273: div <= 91575;
				274: div <= 91241;
				275: div <= 90909;
				276: div <= 90580;
				277: div <= 90253;
				278: div <= 89928;
				279: div <= 89606;
				280: div <= 89286;
				281: div <= 88968;
				282: div <= 88652;
				283: div <= 88339;
				284: div <= 88028;
				285: div <= 87719;
				286: div <= 87413;
				287: div <= 87108;
				288: div <= 86806;
				289: div <= 86505;
				290: div <= 86207;
				291: div <= 85911;
				292: div <= 85616;
				293: div <= 85324;
				294: div <= 85034;
				295: div <= 84746;
				296: div <= 84459;
				297: div <= 84175;
				298: div <= 83893;
				299: div <= 83612;
				300: div <= 83333;
				301: div <= 83056;
				302: div <= 82781;
				303: div <= 82508;
				304: div <= 82237;
				305: div <= 81967;
				306: div <= 81699;
				307: div <= 81433;
				308: div <= 81169;
				309: div <= 80906;
				310: div <= 80645;
				311: div <= 80386;
				312: div <= 80128;
				313: div <= 79872;
				314: div <= 79618;
				315: div <= 79365;
				316: div <= 79114;
				317: div <= 78864;
				318: div <= 78616;
				319: div <= 78370;
				320: div <= 78125;
				512: div <= 48828;
				1024: div <= 24414;
				1200: div <= 20833;
				2048: div <= 12207;
				2400: div <= 10417;
				4096: div <= 6104;
				5120: div <= 4883;
				8192: div <= 3052;
				9600: div <= 2604;
				16384: div <= 1526;
				19200: div <= 1302;
				32768: div <= 763;
				38400: div <= 651;
				57600: div <= 434;
				65536: div <= 381;
				115200: div <= 217;
				131072: div <= 191;
				250000: div <= 100;
				262144: div <= 95;
				500000: div <= 50;
				524288: div <= 48;
				1048576: div <= 24;
				2097152: div <= 12;
				4194304: div <= 6;
				8388608: div <= 3;
				16777216: div <= 1;			
				default: div <= 25000000;
			endcase
		
		if(wait1 >= div) begin // Divider is divided by 2
			wait1 <= 0; // reset clock
			CLK_ <= ~CLK_;
		end
	 end

endmodule
